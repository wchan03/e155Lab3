// Wava Chan
// wchan@g.hmc.edu
// Sept. 15, 2025
// Testing of Lab 3 for E155

`timescale 1ns/1ps

module lab3_wc_testbench();
	
	// set up all necessary logic 
	
	//generate clock
	
	// instantiate DUT 
	
	//run tests
	
endmodule 